-- ************************************************************************* --
-- PCI�^�[�Q�b�g8 (�o�[�X�g�]���Ή�)
-- ************************************************************************* --
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity PCI_TGT8 is
	port(

	-- PCI�o�X�M���s��(�^�[�Q�b�g8�Ŏg�p����M��) --
		PCICLK		: in	std_logic;			-- PCI�o�X�N���b�N
		RST_n		: in	std_logic;			-- �񓯊����Z�b�g
		PCIAD		: inout	std_logic_vector(31 downto 0);	-- �A�h���X/�f�[�^�o�X
		C_BE_n		: in	std_logic_vector(3 downto 0);	-- PCI�o�X�R�}���h/�o�C�g�C�l�[�u��
		FRAME_n		: in	std_logic;			-- �t���[��
		IRDY_n		: in	std_logic;			-- �C�j�V�G�[�^���f�B
		DEVSEL_n	: out	std_logic;			-- �f�o�C�X�Z���N�V����
		TRDY_n		: out	std_logic;			-- �^�[�Q�b�g���f�B
		STOP_n		: out	std_logic;			-- �]���X�g�b�v�v��
		PAR			: inout	std_logic;			-- �p���e�B�r�b�g
		IDSEL		: in	std_logic;			-- �R���t�B�O���[�V�����f�o�C�X�Z���N�g
		INTA_n		: out	std_logic;			-- ���荞�ݏo�� INTA#

	-- PCI�o�X�M���s��(�^�[�Q�b�g8�Ŗ��g�p�ȐM��) --
		PERR_n		: out	std_logic;			-- �p���e�B�G���[
		SERR_n		: out	std_logic;			-- �V�X�e���G���[
		REQ_n		: out	std_logic;			-- �o�X�g�p�v���M��
		GNT_n		: in	std_logic;			-- �o�X�g�p�����M��
		INTB_n		: out	std_logic;			-- ���荞�ݏo�� INTB#
		INTC_n		: out	std_logic;			-- ���荞�ݏo�� INTC#
		INTD_n		: out	std_logic;			-- ���荞�ݏo�� INTD#

	-- ���[�J���o�X�M���s��
		MEM_ADRS	: out	std_logic_vector(23 downto 0);	-- �������A�h���X�o�X
		MEM_DATA	: inout	std_logic_vector(31 downto 0);	-- �������f�[�^�o�X
		MEM_CEn		: out	std_logic;			-- SRAM0�`3 /CE
		MEM_OEn		: out	std_logic;			-- SRAM0�`3 /OE
		MEM_WE0n	: out	std_logic;			-- SRAM0 /WE
		MEM_WE1n	: out	std_logic;			-- SRAM1 /WE
		MEM_WE2n	: out	std_logic;			-- SRAM2 /WE
		MEM_WE3n	: out	std_logic;			-- SRAM3 /WE

	-- �O�����荞�ݓ��̓s��
		INT_IN3		: in	std_logic;			-- ���荞�ݓ���3
		INT_IN2		: in	std_logic;			-- ���荞�ݓ���2
		INT_IN1		: in	std_logic;			-- ���荞�ݓ���1
		INT_IN0		: in	std_logic			-- ���荞�ݓ���0

	);
end entity PCI_TGT8;

architecture RTL of PCI_TGT8 is


-- ************************************************************************* --
-- **********	���W�X�^/�萔 ��`����
-- ************************************************************************* --

-- PCI�o�X�R�}���h/�A�h���X/IDSEL�z�[���h���W�X�^ --
	signal PCI_BusCommand	: std_logic_vector(3 downto 0)		:=	(others => '0');	-- PCI�o�X�R�}���h���W�X�^
	signal PCI_Address	: std_logic_vector(31 downto 0)		:=	(others => '0');	-- PCI�A�h���X���W�X�^
	signal PCI_IDSEL	: std_logic								:=	'0'				;						-- IDSEL���W�X�^

-- ���[�J���o�X�V�[�P���T �X�^�[�g�t���O
	signal LOCAL_Bus_Start : std_logic							:=	'0';
-- ���[�J���o�X�V�[�P���T �f�[�^�]�������t���O
	signal LOCAL_DTACK     : std_logic							:=	'0';

-- �g���C�X�e�[�g�o�b�t�@����p�̃t���b�v�t���b�v��` --
	-- PCI�o�X�M����
	signal PCIAD_HiZ  : std_logic								:=	'1';						-- AD�|�[�g�o�̓h���C�u����
	signal PCIAD_Port : std_logic_vector(31 downto 0)			:=	(others => '0');	-- AD�|�[�g�o�̓��W�X�^
	signal DEVSEL_HiZ, DEVSEL_Port : std_logic					:=	'1';	-- DEVSEL#�o�̓h���C�u����/�o�̓��W�X�^
	signal TRDY_HiZ, TRDY_Port     : std_logic					:=	'1';	-- TRDY#�o�̓h���C�u����/�o�̓��W�X�^
	signal INTA_HiZ                : std_logic					:=	'1';	-- INTA#�o�̓h���C�u����/�o�̓��W�X�^
	signal INTA_Port               : std_logic					:=	'0';	-- INTA#�o�̓h���C�u����/�o�̓��W�X�^
	signal PAR_HiZ                 : std_logic					:=	'1';	-- PAR�o�̓h���C�u����/�o�̓��W�X�^
	signal PAR_Port                : std_logic					:=	'0';	-- PAR�o�̓h���C�u����/�o�̓��W�X�^
	signal STOP_HiZ, STOP_Port     : std_logic					:=	'1';	-- STOP�o�̓h���C�u����/�o�̓��W�X�^
		
		
	--	signal PERR_HiZ, PERR_Port     : std_logic;	-- �_�~�[�m�[�h(�^�[�Q�b�g8���g�p)
	--	signal SERR_HiZ, SERR_Port     : std_logic;
	--	signal REQ_HiZ,  REQ_Port      : std_logic;
	--	signal INTB_HiZ, INTB_Port     : std_logic;
	--	signal INTC_HiZ, INTC_Port     : std_logic;
	--	signal INTD_HiZ, INTD_Port     : std_logic;

--  PCI�o�X�R�}���h(�r�b�g�p�^�[����`) --
	-- �R���t�B�M�����[�V�����T�C�N��
	constant PCI_CfgCycle      : std_logic_vector(3 downto 1) := ("101");
	constant PCI_CfgReadCycle  : std_logic_vector(3 downto 0) := ("1010");
	constant PCI_CfgWriteCycle : std_logic_vector(3 downto 0) := ("1011");
	-- �������T�C�N��
	constant PCI_MemCycle      : std_logic_vector(3 downto 1) := ("011");
	constant PCI_MemReadCycle  : std_logic_vector(3 downto 0) := ("0110");
	constant PCI_MemWriteCycle : std_logic_vector(3 downto 0) := ("0111");
	-- I/O�T�C�N��
	constant PCI_IoCycle       : std_logic_vector(3 downto 1) := ("001");
	constant PCI_IoReadCycle   : std_logic_vector(3 downto 0) := ("0010");
	constant PCI_IoWriteCycle  : std_logic_vector(3 downto 0) := ("0011");

-- �R���t�B�M�����[�V�������W�X�^�Q(�ǂݏo����p���W�X�^) --
--	constant CFG_VendorID   : std_logic_vector(15 downto 0) := (X"6809");	-- �x���_ID   6809h
--	constant CFG_DeviceID   : std_logic_vector(15 downto 0) := (X"8000");	-- �f�o�C�XID 8000h
--	constant CFG_Command    : std_logic_vector(15 downto 0) := (X"0000");
--	constant CFG_Status     : std_logic_vector(15 downto 0) := (X"0200");	-- DEVSEL# ��������
--	constant CFG_BaseClass  : std_logic_vector(7  downto 0) := (X"05");		-- 05h RAM
--	--constant CFG_BaseClass  : std_logic_vector(7  downto 0) := (X"FF");		-- 05h RAM
--	constant CFG_SubClass   : std_logic_vector(7  downto 0) := (X"00");
--	constant CFG_ProgramIF  : std_logic_vector(7  downto 0) := (X"00");
--	constant CFG_RevisionID : std_logic_vector(7  downto 0) := (X"01");		-- ���r�W���� 1
--	constant CFG_HeaderType : std_logic_vector(7  downto 0) := (X"00");		-- �w�b�_�^�C�v0
--	constant CFG_Int_Pin    : std_logic_vector(7  downto 0) := (X"01");		-- INTA#�̂ݎg�p
	
	-- �R���t�B�M�����[�V�������W�X�^�Q(�ǂݏo����p���W�X�^) -- hong pci
	constant CFG_VendorID   : std_logic_vector(15 downto 0) := (X"1172");	-- �x���_ID	
	constant CFG_DeviceID   : std_logic_vector(15 downto 0) := (X"0004");	-- �f�o�C�XID
	constant CFG_Command    : std_logic_vector(15 downto 0) := (X"0000");
	constant CFG_Status     : std_logic_vector(15 downto 0) := (X"0200");	-- DEVSEL# ��������
	constant CFG_BaseClass  : std_logic_vector(7  downto 0) := (X"FF");		-- 05h RAM
	constant CFG_SubClass   : std_logic_vector(7  downto 0) := (X"00");
	constant CFG_ProgramIF  : std_logic_vector(7  downto 0) := (X"00");
	constant CFG_RevisionID : std_logic_vector(7  downto 0) := (X"01");		-- ���r�W���� 1
	constant CFG_HeaderType : std_logic_vector(7  downto 0) := (X"00");		-- �w�b�_�^�C�v0
	constant CFG_Int_Pin    : std_logic_vector(7  downto 0) := (X"01");		-- INTA#�̂ݎg�p
	
	

-- �R���t�B�M�����[�V�������W�X�^�Q(�ǂݏ������W�X�^) --
	-- �R�}���h���W�X�^ �������C�l�[�u���r�b�g
	signal CFG_Cmd_Mem : std_logic						:=	'0';
	-- �R�}���h���W�X�^ I/O�C�l�[�u���r�b�g
	signal CFG_Cmd_Io : std_logic						:=	'0';
	-- �R�}���h���W�X�^ ���荞�݃f�B�Z�[�u���r�b�g
	signal CFG_Cmd_IntDis : std_logic					:=	'0';
	-- �X�e�[�^�X���W�X�^ ���荞�݃X�e�[�^�X�r�b�g
	signal CFG_Sta_IntSta : std_logic					:=	'0';
	-- �x�[�X�A�h���X���W�X�^(���������)
	signal CFG_Base_Addr0 : std_logic_vector(31 downto 24)	:=	(others => '0');
	-- �x�[�X�A�h���X���W�X�^(I/O���)
	signal CFG_Base_Addr1 : std_logic_vector(15 downto 2)		:=	(others => '0');
	-- �C���^���v�g���C�����W�X�^
	signal CFG_Int_Line : std_logic_vector(7 downto 0)	:=	(others => '0');
	
		
		
-- �A�h���X�f�R�[�h�t���O
	signal Hit_Device : std_logic			:=	'0'	;	-- �f�o�C�X�q�b�g
	signal Hit_Memory : std_logic			:=	'0'	;	-- �������T�C�N���q�b�g
	signal Hit_Io : std_logic				:=	'0'	;		-- I/O�T�C�N���q�b�g
	signal Hit_Config : std_logic			:=	'0'	;	-- �R���t�B�O���[�V�����T�C�N���q�b�g

-- PCIAD�o�X�h���C�u���p���e�B�v�Z
	signal TGT_PAR    : std_logic			:=	'0'	;

-- ���[�J���o�X �g���C�X�e�[�g����
	signal MEM_DATA_HiZ  : std_logic		:=	'0'	;	-- �������f�[�^�o�X�g���C�X�e�[�g����
	signal MEM_DATA_Port : std_logic_vector(31 downto 0)	:=	(others => '0');	-- �������f�[�^�o�X

	
		
--  ���荞�ݐ��䃌�W�X�^�Q
	-- ���荞�݃X�e�[�^�X/�t���O���W�X�^
	signal INT_STAT3 : std_logic			:=	'0'	;
	signal INT_STAT2 : std_logic			:=	'0'	;
	signal INT_STAT1 : std_logic			:=	'0'	;
	signal INT_STAT0 : std_logic			:=	'0'	;
	-- ���荞�݃}�X�N(����)���W�X�^
	signal INT_MSK3 : std_logic			:=	'0'	;
	signal INT_MSK2 : std_logic			:=	'0'	;
	signal INT_MSK1 : std_logic			:=	'0'	;
	signal INT_MSK0 : std_logic			:=	'0'	;
	-- ���荞�݃X�e�[�^�X�N���A�w�����W�X�^
	signal INT_CLR3 : std_logic			:=	'0'	;
	signal INT_CLR2 : std_logic			:=	'0'	;
	signal INT_CLR1 : std_logic			:=	'0'	;
	signal INT_CLR0 : std_logic			:=	'0'	;
	
	signal wPCI_CURRENT_STATE	: std_logic_vector (2 downto 0)	:=	(others => '0');	-- ���݂̃X�e�[�g
	
		
begin


-- ************************************************************************* --
-- **********	����������
-- ************************************************************************* --

-- �g���C�X�e�[�g�o�b�t�@����
	MEM_DATA <= (others => 'Z') when MEM_DATA_HiZ = '1' else MEM_DATA_Port;
	PCIAD    <= (others => 'Z') when PCIAD_HiZ = '1'    else PCIAD_Port;
	DEVSEL_n <= 'Z'	when DEVSEL_HiZ = '1'	else DEVSEL_Port;
	TRDY_n   <= 'Z'	when TRDY_HiZ = '1'	else TRDY_Port;
	INTA_n <= 'Z'	when INTA_HiZ = '1'	else INTA_Port; INTA_Port <= '0';
	PAR    <= 'Z'	when PAR_HiZ  = '1'	else PAR_Port;
	STOP_n <= 'Z'	when STOP_HiZ = '1'	else STOP_Port;

-- ���g�p�s���̏�Ԑݒ�(�n�C�C���s�[�_���X��ԂɌŒ�)
	PERR_n <= 'Z'		;	--	when PERR_HiZ = '1'	else PERR_Port; PERR_HiZ <= '1'; PERR_Port <= '0';
	SERR_n <= 'Z'		;	--	when SERR_HiZ = '1'	else SERR_Port; SERR_HiZ <= '1'; SERR_Port <= '0';
	REQ_n  <= 'Z'		;	--	when REQ_HiZ  = '1'	else REQ_Port;	REQ_HiZ  <= '0'; REQ_Port  <= '1';
	INTB_n <= 'Z'		;	--	when INTB_HiZ = '1'	else INTB_Port; INTB_HiZ <= '1'; INTB_Port <= '0';
	INTC_n <= 'Z'		;	--	when INTC_HiZ = '1'	else INTC_Port; INTC_HiZ <= '1'; INTC_Port <= '0';
	INTD_n <= 'Z'		;	--	when INTD_HiZ = '1'	else INTD_Port; INTD_HiZ <= '1'; INTD_Port <= '0';
	
-- ************************************************************************* --
-- **********	PCI�^�[�Q�b�g�V�[�P���T
-- ************************************************************************* --

PCI_TGT_Seq : process( PCICLK, RST_n )

-- PCI�^�[�Q�b�g�V�[�P���T �X�e�[�g�o�����[���W�X�^ --
	variable PCI_CURRENT_STATE	: std_logic_vector (2 downto 0)		:=	(others => '0')	;	-- ���݂̃X�e�[�g
	variable PCI_NEXT_STATE		: std_logic_vector (2 downto 0)	:=	(others => '0')	;	-- ���̃X�e�[�g

-- PCI�^�[�Q�b�g�V�[�P���T �X�e�[�g�}�V����`
	constant BUS_IDLE		: std_logic_vector (2 downto 0) :="000";
	constant ADRS_COMPARE	: std_logic_vector (2 downto 0) :="001";
	constant BUS_BUSY		: std_logic_vector (2 downto 0) :="010";
	constant WAIT_IRDY		: std_logic_vector (2 downto 0) :="011";
	constant WAIT_LOCAL_ACK : std_logic_vector (2 downto 0) :="100";
	constant ACC_COMPLETE	: std_logic_vector (2 downto 0) :="101";
	constant DIS_CONNECT	: std_logic_vector (2 downto 0) :="110";
	constant TURN_AROUND	: std_logic_vector (2 downto 0) :="111";

begin

-- ********** ���Z�b�g������ ********** --
	if (RST_n = '0') then	-- PCI�o�X���Z�b�g��(�񓯊����Z�b�g)

		PCI_CURRENT_STATE	:= BUS_IDLE;	-- �X�e�[�g�}�V�� IDLE��� ���Z�b�g
		PCI_NEXT_STATE		:= BUS_IDLE;	-- �X�e�[�g�}�V�� IDLE��� ���Z�b�g

		LOCAL_Bus_Start <= '0';		-- ���[�J���o�X�V�[�P���T �X�^�[�g�t���O �N���A

		PCI_BusCommand <= (others => '0');	-- PCI�o�X�R�}���h���W�X�^ �N���A
		PCI_Address <= (others => '0');		-- PCI�o�X�A�h���X���W�X�^ �N���A
		PCI_IDSEL <= '0';					-- IDSEL���W�X�^ �N���A

	-- ����o�͒[�q���n�C�C���s�[�_���X
		PCIAD_HiZ <= '1';
		DEVSEL_HiZ <= '1'; DEVSEL_Port <= '1';	-- DEVSEL#="H"
		TRDY_HiZ   <= '1'; TRDY_Port   <= '1';	-- TRDY#="H"
		STOP_HiZ   <= '1'; STOP_Port   <= '1';	-- STOP#="H"


-- ********** PCI�^�[�Q�b�g�V�[�P���T �X�e�[�g�}�V�� ********** --
	elsif (PCICLK'event and PCICLK = '1') then

		PCI_CURRENT_STATE := PCI_NEXT_STATE;	-- �X�e�[�g�}�V������
		case PCI_CURRENT_STATE is

	-- ********** BUS_IDLE���̓��� ********** --
		when BUS_IDLE =>	-- �g�����U�N�V�����̊J�n�҂�

			if (FRAME_n = '0' and IRDY_n /= '0') then	-- �g�����U�N�V�����J�n
				PCI_BusCommand <= C_BE_n;	-- PCI�o�X�R�}���h�擾
				PCI_Address <= PCIAD;		-- �A�h���X�擾
				PCI_IDSEL <= IDSEL;			-- IDSEL�擾
				PCI_NEXT_STATE := ADRS_COMPARE;

			else	-- �o�X�A�C�h�������̃X�e�[�g�ɂƂǂ܂�
				PCI_NEXT_STATE := BUS_IDLE;
			end if;


	-- ********** ADRS_COMPARE���̓��� ********** --
		when ADRS_COMPARE =>	-- �A�h���X�f�R�[�h���ʂ𒲂ׂ�

			if (Hit_Device = '1') then	-- �������I�����ꂽ
				DEVSEL_Port <= '0'; DEVSEL_HiZ <= '0';	-- DEVLSEL#�A�T�[�g
				TRDY_HiZ <= '0';	-- TRDY# �� "H"�Ƀh���C�u
				STOP_HiZ <= '0';	-- STOP# �� "H"�Ƀh���C�u
				PCI_NEXT_STATE := WAIT_IRDY;	-- �C�j�V�G�[�^���f�B��҂X�e�[�g��

			else	-- �������I������Ă��Ȃ�
				PCI_NEXT_STATE := BUS_BUSY;	-- �g�����U�N�V�����̏I����҂X�e�[�g��
			end if;


	-- ********** BUS_BUSY���̓��� ********** --
		when BUS_BUSY =>	-- �g�����U�N�V�����I���҂�

			if (FRAME_n = '1' and IRDY_n = '1') then	-- �g�����U�N�V�����I��(�A�C�h��)
				PCI_NEXT_STATE := BUS_IDLE;	-- �g�����U�N�V�����J�n�҂��X�e�[�g��

			else	-- �g�����U�N�V�������Ȃ炱�̃X�e�[�g�ɂƂǂ܂�
				PCI_NEXT_STATE := BUS_BUSY;
			end if;


	-- ********** WAIT_IRDY���̓��� ********** --
		when WAIT_IRDY =>	-- �C�j�V�G�[�^���f�B�҂�

			if (IRDY_n = '0') then	-- �C�j�V�G�[�^�̏�������
				if (PCI_BusCommand(0) = '0') then	-- ���[�h�T�C�N���̂Ƃ�
					PCIAD_HiZ <= '0' ;				-- PCIAD[31:0]�o�X�h���C�u
				end if;
				LOCAL_Bus_Start <= '1';	-- ���[�J���o�X�V�[�P���T �X�^�[�g!
				PCI_NEXT_STATE := WAIT_LOCAL_ACK;	-- ���[�J���o�X�V�[�P���T�I���҂��X�e�[�g��

			else	-- �C�j�V�G�[�^�̏������܂��Ȃ炱�̃X�e�[�g�ɂƂǂ܂�
				PCI_NEXT_STATE := WAIT_IRDY;
			end if;


	-- ********** WAIT_LOCAL_ACK���̓��� ********** --
		when WAIT_LOCAL_ACK =>	-- ���[�J���o�X�V�[�P���T�I���҂�

			LOCAL_Bus_Start <= '0';	-- ���[�J���o�X�V�[�P���T �X�^�[�g�t���O �N���A

			if (LOCAL_DTACK = '1') then	-- ���[�J���o�X�V�[�P���T �f�[�^�]������
				TRDY_Port <= '0';	-- TRDY# �A�T�[�g
				PCI_NEXT_STATE := ACC_COMPLETE;	-- �A�N�Z�X�����X�e�[�g��

			else	-- ���[�J���o�X�V�[�P���T�̏������܂��Ȃ炱�̃X�e�[�g�ɂƂǂ܂�
				PCI_NEXT_STATE := WAIT_LOCAL_ACK;
			end if;


	-- ********** ACC_COMPLETE���̓��� ********** --
		when ACC_COMPLETE =>	-- �A�N�Z�X�����X�e�[�g

			TRDY_Port <= '1';		-- TRDY# �f�B�A�T�[�g
			PCIAD_HiZ <= '1' ;		-- PCIAD[31:0]�o�X�h���C�u���

			if (FRAME_n = '0') then			-- FRAME# = 'L'�Ȃ�o�[�X�g�]���v��

				if ( Hit_Memory = '1' and PCI_Address(1 downto 0) = "00"
						-- ���������&�A�h���X�C���N�������g���[�h=���j�A�o�[�X�g
						-- �o�[�X�g�]���A�h���X���ŏ�ʈȊO�Ȃ�
						and PCI_Address(23 downto 2) /= "1111111111111111111111") then
									-- �A�h���X���ŏI�A�h���X�ł͂Ȃ�
					PCI_Address(23 downto 2) <= PCI_Address(23 downto 2) + '1';
					PCI_NEXT_STATE := WAIT_IRDY;	-- �C�j�V�G�[�^���f�B��҂X�e�[�g��

				else
					STOP_Port <= '0';	-- STOP# �A�T�[�g
					PCI_NEXT_STATE := DIS_CONNECT;	-- �f�B�X�R�l�N�g�X�e�[�g��
				end if;

			else	-- �P��f�[�^�t�F�[�Y�̃g�����U�N�V�����̎�
				DEVSEL_Port <= '1';		-- DEVSEL#�f�B�A�T�[�g
				PCI_NEXT_STATE := TURN_AROUND;	--  �^�[���A���E���h�X�e�[�g��
			end if;


	-- ********** DIS_CONNECT���̓��� ********** --
		when DIS_CONNECT =>		-- �f�B�X�R�l�N�g����

			if (FRAME_n = '1') then	-- �C�j�V�G�[�^��STOP#��F��
				DEVSEL_Port <= '1';	-- DEVSEL# �f�B�A�T�[�g
				STOP_Port <= '1';	-- STOP# �f�B�A�T�[�g
				PCI_NEXT_STATE := TURN_AROUND;	-- ����TURN_AROUND�X�e�[�g��

			else	-- �C�j�V�G�[�^��STOP#��F�����Ă��Ȃ���΂��̃X�e�[�g�ɂƂǂ܂�
				PCI_NEXT_STATE := DIS_CONNECT;
			end if;


	-- ********** TURN_AROUND���̓��� ********** --
		when TURN_AROUND =>		-- �^�[���A���E���h�X�e�[�g

			DEVSEL_HiZ <= '1';			-- DEVSEL#�h���C�u���
			TRDY_HiZ <= '1';			-- TRDY#�h���C�u���
			STOP_HiZ <= '1';			-- STOP#�h���C�u���
			PCI_NEXT_STATE := BUS_IDLE;	-- �g�����U�N�V�����J�n�҂��X�e�[�g��


	-- ****************************************** --
		when others => null;	-- ����ȊO�̒l�ł͉������Ȃ��ꍇ�ł��K�������

	end case;

	end if;

	wPCI_CURRENT_STATE	<=	PCI_CURRENT_STATE	;
	
end process PCI_TGT_Seq;



-- ************************************************************************* --
-- **********	���[�J���o�X�V�[�P���T
-- ************************************************************************* --
MEM_ADRS(23 downto 2) <= PCI_Address(23 downto 2);
MEM_ADRS(1 downto 0) <=	"00";
LOCAL_BUS_Seq : process(PCICLK, RST_n)

-- ���[�J���o�X�V�[�P���T �X�e�[�g�o�����[���W�X�^ --
	variable LOCAL_CURRENT_STATE : std_logic_vector (2 downto 0)	:= (others => '0')	;	-- ���݂̃X�e�[�g
	variable LOCAL_NEXT_STATE : std_logic_vector (2 downto 0)	:= (others => '0')	;		-- ���̃X�e�[�g

-- ���[�J���o�X�V�[�P���T �X�e�[�g�}�V����`
	constant LOCAL_IDLE			: std_logic_vector(2 downto 0) := "000";
	constant LOCAL_MEM_ACCESS	: std_logic_vector(2 downto 0) := "001";
	constant LOCAL_IO_ACCESS	: std_logic_vector(2 downto 0) := "010";
	constant LOCAL_CFG_ACCESS	: std_logic_vector(2 downto 0) := "011";
	constant LOCAL_STATE_COMP	: std_logic_vector(2 downto 0) := "100";

-- �������A�N�Z�X �E�F�C�g�J�E���^
	variable WAIT_Count : std_logic_vector(3 downto 0)		:=	(others => '0');

begin

-- ********** ���Z�b�g������ ********** --
	if (RST_n = '0') then	-- PCI�o�X���Z�b�g���A�T�[�g���ꂽ�Ƃ�

		-- �X�e�[�g�o�����[���W�X�^�N���A
		LOCAL_CURRENT_STATE := (others => '0');	-- ���[�J���o�X�V�[�P���T ���Z�b�g
		LOCAL_NEXT_STATE := (others => '0');	-- ���[�J���o�X�V�[�P���T ���Z�b�g

		-- �R���t�B�O���[�V�������W�X�^ ���[�h/���C�g���W�X�^ �C���^���v�g���C�� �N���A
		CFG_Cmd_Mem <= '0';
		CFG_Cmd_Io  <= '0';
		CFG_Cmd_IntDis <= '0';
		CFG_Base_Addr0 <= (others => '0');
		CFG_Base_Addr1 <= (others => '0');
		CFG_Int_Line <= (others => '0');

		-- ���[�J���o�X������f�B�Z�[�u��
		MEM_CEn  <= '1';	-- SRAM0�`3 /CE
		MEM_OEn  <= '1';	-- SRAM0�`3 /OE
		MEM_WE0n <= '1';	-- SRAM0 /WE
		MEM_WE1n <= '1';	-- SRAM1 /WE
		MEM_WE2n <= '1';	-- SRAM2 /WE
		MEM_WE3n <= '1';	-- SRAM3 /WE
		MEM_DATA_HiZ  <= '0';	-- �f�[�^�o�X�o�͕���

		PCIAD_Port <= (others => '0');		-- AD�o�̓��W�X�^ �N���A
		MEM_DATA_Port <= (others => '0');	-- MEM_DATA�o�̓��W�X�^ �N���A

		-- �������A�N�Z�X �E�F�C�g�J�E���^ �N���A
		WAIT_Count := (others => '0');

		-- ���[�J���o�X�V�[�P���T �f�[�^�]�������t���O �N���A
		LOCAL_DTACK <= '0';

		-- ���荞�ݐ��䃌�W�X�^ --
		INT_MSK3 <= '0';	-- ���荞�݃}�X�N���W�X�^ �N���A
		INT_MSK2 <= '0';
		INT_MSK1 <= '0';
		INT_MSK0 <= '0';
		INT_CLR3 <= '0';	-- ���荞�݃X�e�[�^�X�N���A�w���M�� �N���A
		INT_CLR2 <= '0';
		INT_CLR1 <= '0';
		INT_CLR0 <= '0';


-- ********** ���[�J���o�X�V�[�P���T �X�e�[�g�}�V�� ********** --
	elsif (PCICLK'event and PCICLK = '1') then

		LOCAL_CURRENT_STATE := LOCAL_NEXT_STATE;
		case LOCAL_CURRENT_STATE is

	-- ********** LOCAL_IDLE���̓��� ********** --
		when LOCAL_IDLE =>	-- ���[�J���o�X�V�[�P���T �X�^�[�g�w���҂�

			if (LOCAL_Bus_Start = '1' ) then	-- ���[�J���o�X�V�[�P���T �X�^�[�g!

				if (Hit_Config = '1') then	-- �R���t�B�O���[�V�����T�C�N���q�b�g
					LOCAL_NEXT_STATE := LOCAL_CFG_ACCESS;	-- �R���t�B�O���[�V�����X�e�[�g��
				end if;
				if (Hit_Memory = '1') then	-- �������T�C�N���q�b�g
					LOCAL_NEXT_STATE := LOCAL_MEM_ACCESS;	-- �������A�N�Z�X�X�e�[�g��
				end if;
				if (Hit_Io = '1') then		-- I/O�T�C�N���q�b�g
					LOCAL_NEXT_STATE := LOCAL_IO_ACCESS;	-- I/O�A�N�Z�X�X�e�[�g��
				end if;

			else	-- ���[�J���o�X�V�[�P���T �X�^�[�g�t���O���܂��Ȃ炱�̃X�e�[�g�ɂƂǂ܂�

				LOCAL_NEXT_STATE := LOCAL_IDLE;
			end if;


	-- ********** LOCAL_MEM_ACCESS���̓��� ********** --
		when LOCAL_MEM_ACCESS =>

			case WAIT_Count is
			when X"0" =>	-- �E�F�C�g�J�E���^0�N���b�N��
				MEM_CEn <= '0';		-- SRAM /CE �A�T�[�g
				if (PCI_BusCommand(0) = '1') then	-- ���������C�g�T�C�N��
					MEM_DATA_Port(31 downto 0) <= PCIAD(31 downto 0); -- ���C�g�f�[�^
				else						-- ���������[�h�T�C�N��
					MEM_DATA_HiZ <= '1';	-- ���[�J���f�[�^�o�X���͕���
				end if;
				LOCAL_NEXT_STATE := LOCAL_MEM_ACCESS;	-- �������A�N�Z�X�͂܂��I���Ȃ�

			when X"1" =>	-- �E�F�C�g�J�E���^1�N���b�N��
				if (PCI_BusCommand(0) = '1') then	-- ���������C�g�T�C�N��
					MEM_WE3n <= C_BE_n(3);	-- �o�C�g�C�l�[�u����/WE�ɏo��
					MEM_WE2n <= C_BE_n(2);
					MEM_WE1n <= C_BE_n(1);
					MEM_WE0n <= C_BE_n(0);
				else						-- ���������[�h�T�C�N��
					MEM_OEn <= '0';			-- SRAM /OE �A�T�[�g
				end if;
				LOCAL_NEXT_STATE := LOCAL_MEM_ACCESS;	-- �������A�N�Z�X�͂܂��I���Ȃ�

			when X"4" =>	-- �E�F�C�g�J�E���^4�N���b�N��
				if (PCI_BusCommand(0) = '1') then	-- ���������C�g�T�C�N��
					MEM_WE3n <= '1';	-- SRAM /WE �f�B�Z�[�u��
					MEM_WE2n <= '1';
					MEM_WE1n <= '1';
					MEM_WE0n <= '1';
				else									-- ���������[�h�T�C�N��
					PCIAD_Port(31 downto 0) <= MEM_DATA;-- SRAM�f�[�^��AD�o�X�ɏo��
					MEM_OEn <= '1';						-- SRAM /OE �f�B�A�T�[�g
				end if;
				LOCAL_DTACK <= '1';		-- ���[�J���o�X�V�[�P���T �f�[�^�]�������t���O �Z�b�g
				LOCAL_NEXT_STATE := LOCAL_STATE_COMP;	-- �������A�N�Z�X����

			when others =>	-- ���̂܂܂̏�ԂŃE�F�C�g���Ԃ��o�߂���̂�҂�
				LOCAL_NEXT_STATE := LOCAL_MEM_ACCESS;	-- �������A�N�Z�X�͂܂��I���Ȃ�

			end case;

			WAIT_Count := WAIT_Count + '1';	-- �E�F�C�g�J�E���g + 1


		-- ********** LOCAL_IO_ACCESS���̓��� ********** --
		when LOCAL_IO_ACCESS =>

			if (PCI_BusCommand(0) = '1') then	-- ���C�g�T�C�N��

				case PCI_Address(1 downto 0) is
					when "00" =>				-- ���荞�݃X�e�[�^�X���W�X�^�ւ̃A�N�Z�X
						INT_CLR3 <= PCIAD(3);		-- �X�e�[�^�X�N���A #3
						INT_CLR2 <= PCIAD(2);		-- �X�e�[�^�X�N���A #2
						INT_CLR1 <= PCIAD(1);		-- �X�e�[�^�X�N���A #1
						INT_CLR0 <= PCIAD(0);		-- �X�e�[�^�X�N���A #0

					when "10" =>				-- ���荞�݃}�X�N���W�X�^�ւ̃A�N�Z�X
						INT_MSK3 <= PCIAD(19);		-- ���荞�݃}�X�N #3
						INT_MSK2 <= PCIAD(18);		-- ���荞�݃}�X�N #2
						INT_MSK1 <= PCIAD(17);		-- ���荞�݃}�X�N #1
						INT_MSK0 <= PCIAD(16);		-- ���荞�݃}�X�N #0

					when others => null;		-- ����ȊO�̃A�N�Z�X�͖���
				end case;

			else	-- ���[�h�T�C�N��

				case PCI_Address(1 downto 0) is
					when "00" =>				-- ���荞�݃X�e�[�^�X���W�X�^�ւ̃A�N�Z�X
						PCIAD_Port(31 downto  4) <= (others => '0');
						PCIAD_Port(3)  <= INT_STAT3;-- ���荞��3�X�e�[�^�X
						PCIAD_Port(2)  <= INT_STAT2;-- ���荞��2�X�e�[�^�X
						PCIAD_Port(1)  <= INT_STAT1;-- ���荞��1�X�e�[�^�X
						PCIAD_Port(0)  <= INT_STAT0;-- ���荞��0�X�e�[�^�X

					when "10" =>				-- ���荞�݃}�X�N���W�X�^�ւ̃A�N�Z�X
						PCIAD_Port(31 downto 20) <= (others => '0');
						PCIAD_Port(19) <= INT_MSK3;	-- ���荞��3�}�X�N
						PCIAD_Port(18) <= INT_MSK2;	-- ���荞��2�}�X�N
						PCIAD_Port(17) <= INT_MSK1;	-- ���荞��1�}�X�N
						PCIAD_Port(16) <= INT_MSK0;	-- ���荞��0�}�X�N
						PCIAD_Port(15 downto  4) <= (others => '0');

					when others =>				-- ����ȊO�̃A�N�Z�X��0��Ԃ�
						PCIAD_Port(31 downto 0) <= (others => '0');
				end case;

			end if;

			LOCAL_DTACK <= '1';
			LOCAL_NEXT_STATE := LOCAL_STATE_COMP;


	-- ********** LOCAL_CFG_ACCESS���̓��� ********** --
		when LOCAL_CFG_ACCESS =>	-- �R���t�B�O���[�V�����T�C�N��

			if (PCI_BusCommand(0) = '1' ) then	-- �R���t�B�O���[�V�������C�g�T�C�N��

				case PCI_Address(7 downto 2) is

				when "000001" =>	-- �R�}���h���W�X�^
					if (C_BE_n(1) = '0') then
						CFG_Cmd_IntDis <= PCIAD(10);-- ���荞�݃f�B�Z�[�u��
					end if;
					if (C_BE_n(0) = '0') then
						CFG_Cmd_Mem <= PCIAD(1);	-- �������C�l�[�u��
						CFG_Cmd_Io  <= PCIAD(0);	-- I/O�C�l�[�u��
					end if;

				when "000100" =>	-- �x�[�X�A�h���X���W�X�^0
					if (C_BE_n(3) = '0') then
						CFG_Base_Addr0(31 downto 24) <= PCIAD(31 downto 24);
					end if;

				when "000101" =>	-- �x�[�X�A�h���X���W�X�^1
					if (C_BE_n(1) = '0') then
						CFG_Base_Addr1(15 downto  8) <= PCIAD(15 downto  8);
					end if;
					if (C_BE_n(0) = '0') then
						CFG_Base_Addr1( 7 downto  2) <= PCIAD( 7 downto  2);
					end if;

				when "001111" =>	-- ���荞�݃��C�����W�X�^
					if (C_BE_n(0) = '0') then
						CFG_Int_Line(7 downto 0) <= PCIAD(7 downto 0);
					end if;

				when others => null;	-- ����ȊO�̒l�ł͉������Ȃ��ꍇ�ł��K�������

				end case;


			else	-- �R���t�B�O���[�V�������[�h�T�C�N��

				case PCI_Address(7 downto 2) is

				when "000000" =>	-- �x���_ID/�f�o�C�XID
					PCIAD_Port(31 downto 16) <= CFG_DeviceID;
					PCIAD_Port(15 downto  0) <= CFG_VendorID;

				when "000001" =>	-- �R�}���h/�X�e�[�^�X���W�X�^
					PCIAD_Port(31 downto 20) <= CFG_Status(15 downto  4);
					PCIAD_Port(19)           <= CFG_Sta_IntSta;
					PCIAD_Port(18 downto 16) <= CFG_Status( 2 downto  0);
					PCIAD_Port(15 downto 11) <= CFG_Command(15 downto 11);
					PCIAD_Port(10)           <= CFG_Cmd_IntDis;
					PCIAD_Port( 9 downto  2) <= CFG_Command( 9 downto  2);
					PCIAD_Port(1)            <= CFG_Cmd_Mem;
					PCIAD_Port(0)            <= CFG_Cmd_Io;

				when "000010" =>	-- �N���X�R�[�h
					PCIAD_Port(31 downto 24) <= CFG_BaseClass;
					PCIAD_Port(23 downto 16) <= CFG_SubClass;
					PCIAD_Port(15 downto  8) <= CFG_ProgramIF;
					PCIAD_Port( 7 downto  0) <= CFG_RevisionID;

				when "000011" =>	-- �w�b�_�^�C�v�ق�
					PCIAD_Port(31 downto 24) <= (others => '0');
					PCIAD_Port(23 downto 16) <= CFG_HeaderType;
					PCIAD_Port(15 downto  0) <= (others => '0');

				when "000100" =>	-- �x�[�X�A�h���X���W�X�^0
					PCIAD_Port(31 downto 24) <= CFG_Base_Addr0;
					PCIAD_Port(23 downto  0) <= (others => '0');

				when "000101" =>	-- �x�[�X�A�h���X���W�X�^1
					PCIAD_Port(31 downto 16) <= (others => '0');
					PCIAD_Port(15 downto  2) <= CFG_Base_Addr1;
					PCIAD_Port( 1 downto  0) <= "01";

				when "001011" =>	-- �T�u�V�X�e���x���_ID/�T�u�V�X�e��ID
					PCIAD_Port(31 downto 16) <= CFG_DeviceID;
					PCIAD_Port(15 downto  0) <= CFG_VendorID;

				when "001111" =>	-- ���荞�݊֘A���W�X�^
					PCIAD_Port(31 downto 16) <= (others => '0');
					PCIAD_Port(15 downto  8) <= CFG_Int_Pin;
					PCIAD_Port( 7 downto  0) <= CFG_Int_Line;

				when others => -- ���̑��̃��W�X�^
					PCIAD_Port <= (others => '0');	-- ���ׂ�0��Ԃ�

				end case;

			end if;

			LOCAL_DTACK <= '1';		-- ���[�J���o�X�V�[�P���T �f�[�^�]�������t���O �Z�b�g
			LOCAL_NEXT_STATE := LOCAL_STATE_COMP;


	-- ********** LOCAL_STATE_COMP���̓��� ********** --
		when LOCAL_STATE_COMP =>	-- ���[�J���o�X�A�N�Z�X����

			INT_CLR3 <= '0';		-- ���荞�݃N���A�w���M���N���A
			INT_CLR2 <= '0';
			INT_CLR1 <= '0';
			INT_CLR0 <= '0';

			MEM_CEn <= '1';			-- SRAM /CE �f�B�A�T�[�g
			MEM_DATA_HiZ <= '0';	-- ���[�J���f�[�^�o�X�o�͕���
			WAIT_Count := (others => '0');
			LOCAL_DTACK <= '0';		-- ���[�J���o�X�V�[�P���T �f�[�^�]�������t���O �N���A
			LOCAL_NEXT_STATE := LOCAL_IDLE;


	-- ********************************************** --
		when others => null;	-- ����ȊO�̒l�ł͉������Ȃ��ꍇ�ł��K�������

		end case;

	end if;

end process LOCAL_BUS_Seq;



-- ************************************************************************* --
-- **********	���荞�݃R���g���[��
-- ************************************************************************* --

INT_Ctrl : process(PCICLK, RST_n)
	variable INT_IN3_flg1 : std_logic		:=	'0'	;	-- ���荞�ݓ��͏�ԕۑ��t���O
	variable INT_IN2_flg1 : std_logic		:=	'0'	;
	variable INT_IN1_flg1 : std_logic		:=	'0'	;
	variable INT_IN0_flg1 : std_logic		:=	'0'	;
	variable INT_IN3_flg0 : std_logic		:=	'0'	;	-- ���荞�ݓ��͏�ԕۑ��t���O
	variable INT_IN2_flg0 : std_logic		:=	'0'	;
	variable INT_IN1_flg0 : std_logic		:=	'0'	;
	variable INT_IN0_flg0 : std_logic		:=	'0'	;
begin
	if (RST_n = '0') then	-- PCI�o�X���Z�b�g���A�T�[�g���ꂽ�Ƃ�

		INTA_HiZ  <='1';	-- INTA# �n�C�C���s�[�_���X
		CFG_Sta_IntSta <= '0';

		INT_STAT3 <= '0';	-- ���荞�ݗv�����W�X�^ �N���A
		INT_STAT2 <= '0';
		INT_STAT1 <= '0';
		INT_STAT0 <= '0';
		INT_IN3_flg1 := '0';	-- ���荞�ݓ��̓t���O �N���A
		INT_IN2_flg1 := '0';
		INT_IN1_flg1 := '0';
		INT_IN0_flg1 := '0';
		INT_IN3_flg0 := '0';
		INT_IN2_flg0 := '0';
		INT_IN1_flg0 := '0';
		INT_IN0_flg0 := '0';

	elsif (PCICLK'event and PCICLK = '1') then

	-- **********	���荞�݃R���g���[��	 ********** --
		if (INT_CLR3 = '1') then
			INT_STAT3  <= '0';	-- ���荞�݃X�e�[�^�X���W�X�^3�N���A
		elsif (INT_IN3_flg1 = '1' and INT_IN3_flg0 = '0') then	-- �O�����荞�ݓ���3 ��������G�b�W
			INT_STAT3  <= '1';	-- ���荞�݃X�e�[�^�X���W�X�^3
		end if;
		if (INT_CLR2 = '1') then
			INT_STAT2  <= '0';	-- ���荞�݃X�e�[�^�X���W�X�^2�N���A
		elsif (INT_IN2_flg1 = '1' and INT_IN2_flg0 = '0') then	-- �O�����荞�ݓ���2 ��������G�b�W
			INT_STAT2  <= '1';	-- ���荞�݃X�e�[�^�X���W�X�^2
		end if;
		if (INT_CLR1 = '1') then
			INT_STAT1  <= '0';	-- ���荞�݃X�e�[�^�X���W�X�^1�N���A
		elsif (INT_IN1_flg1 = '1' and INT_IN1_flg0 = '0') then	-- �O�����荞�ݓ���1 ��������G�b�W
			INT_STAT1  <= '1';	-- ���荞�݃X�e�[�^�X���W�X�^1
		end if;
		if (INT_CLR0 = '1') then
			INT_STAT0  <= '0';	-- ���荞�݃X�e�[�^�X���W�X�^0�N���A
		elsif (INT_IN0_flg1 = '1' and INT_IN0_flg0 = '0') then	-- �O�����荞�ݓ���0 ��������G�b�W
			INT_STAT0  <= '1';	-- ���荞�݃X�e�[�^�X���W�X�^0
		end if;

		if (
			(CFG_Cmd_IntDis = '0')	-- ���荞�݃f�B�Z�[�u���r�b�g���Z�b�g����Ă��Ȃ�
		) and (
			(INT_STAT3 = '1' and INT_MSK3 = '1') -- �`���l��3���荞�ݔ���&���荞�݉�
			or
			(INT_STAT2 = '1' and INT_MSK2 = '1') -- �`���l��2���荞�ݔ���&���荞�݉�
			or
			(INT_STAT1 = '1' and INT_MSK1 = '1') -- �`���l��1���荞�ݔ���&���荞�݉�
			or
			(INT_STAT0 = '1' and INT_MSK0 = '1') -- �`���l��0���荞�ݔ���&���荞�݉�
		) then
			INTA_HiZ <= '0';	-- INTA#�h���C�u�J�n(�A�T�[�g)
			CFG_Sta_IntSta <= '1';	-- ���荞�ݏo�͒�
		else
			INTA_HiZ <= '1';	-- �n�C�C���s�[�_���X���
			CFG_Sta_IntSta <= '0';
		end if;

		INT_IN3_flg1 := INT_IN3_flg0;
		INT_IN2_flg1 := INT_IN2_flg0;
		INT_IN1_flg1 := INT_IN1_flg0;
		INT_IN0_flg1 := INT_IN0_flg0;
		INT_IN3_flg0 := INT_IN3;	-- ���݂̊��荞�ݓ��͏�Ԃ̕ۑ�
		INT_IN2_flg0 := INT_IN2;
		INT_IN1_flg0 := INT_IN1;
		INT_IN0_flg0 := INT_IN0;

	end if;

end process INT_Ctrl;





-- ************************************************************************* --
-- **********	�A�h���X�f�R�[�_
-- ************************************************************************* --

-- �������T�C�N��or�R���t�B�O���[�V�����T�C�N���q�b�g = �������I������Ă���
Hit_Device <= Hit_Memory or Hit_Config or Hit_Io;

Address_Decoder : process (
				PCI_IDSEL,		-- �R���t�B�O���[�V�����f�o�C�X�Z���N�g
				PCI_Address,	-- PCI�o�X�A�h���X
				PCI_BusCommand,	-- �o�X�R�}���h
				CFG_Base_Addr0,	-- �x�[�X�A�h���X���W�X�^0
				CFG_Base_Addr1,	-- �x�[�X�A�h���X���W�X�^1
				CFG_Cmd_Mem,	-- �R���t�B�O���[�V�������W�X�^ �������C�l�[�u���r�b�g
				CFG_Cmd_Io		-- �R���t�B�O���[�V�������W�X�^ I/O�C�l�[�u���r�b�g
				)
begin

	-- ��������Ԃւ̃A�N�Z�X�A�h���X�ƃx�[�X�A�h���X0����v������
	if (
			PCI_BusCommand(3 downto 1) = PCI_MemCycle	-- �������T�C�N��
		) and (
			PCI_Address(31 downto 24) = CFG_Base_Addr0	-- �x�[�X�A�h���X0�Ɣ�r
		) and (
			CFG_Cmd_Mem = '1'	-- �R���t�B�O���[�V���� �R�}���h���W�X�^ �������C�l�[�u���r�b�g
		)
	then
		Hit_Memory <= '1';	-- �������T�C�N���q�b�g
	else
		Hit_Memory <= '0';
	end if;

	-- I/O��Ԃւ̃A�N�Z�X�A�h���X�ƃx�[�X�A�h���X1����v������
	if (
			PCI_BusCommand(3 downto 1) = PCI_IoCycle	-- I/O�T�C�N��
		) and (
			CFG_Cmd_Io = '1' -- �R���t�B�O���[�V���� �R�}���h���W�X�^ I/O�C�l�[�u���r�b�g
		) and (
			PCI_Address(31 downto 16) = X"0000"		-- ���16�r�b�g��0��
		) and (
			PCI_Address(15 downto 2 ) = CFG_Base_Addr1(15 downto 2)
		)
	then
		Hit_Io <= '1';	-- I/O�T�C�N���q�b�g
	else
		Hit_Io <= '0';
	end if;

	-- �R���t�B�O���[�V������Ԃւ̃A�N�Z�X���ǂ�����F��
	if (
			PCI_BusCommand(3 downto 1) = PCI_CfgCycle	-- �R���t�B�O���[�V�����T�C�N��
		) and (
			PCI_IDSEL = '1'		-- �������I������Ă��邩
		) and (
			PCI_Address(10 downto 8) = "000"	-- �t�@���N�V�����ԍ�0�̂�
		) and (
			PCI_Address(1 downto 0) = "00"		-- �^�C�v0�̂�
		)
	then
		Hit_Config <= '1';	-- �R���t�B�O���[�V�����T�C�N���q�b�g
	else
		Hit_Config <= '0';
	end if;

end process Address_Decoder;



-- ************************************************************************* --
-- **********	�p���e�B�W�F�l���[�^
-- ************************************************************************* --

-- ***** �p���e�B���� ***** --
PCI_Parity_Gen : process (PCIAD_Port, C_BE_n)
	variable temp : std_logic		:=	'0';	-- �e���|����
begin
	-- �^�[�Q�b�g �p���e�B���� --
	temp := '0';
	for I in 0 to 31 loop
		temp := temp xor PCIAD_Port(I);
	end loop;
	TGT_PAR <= temp xor C_BE_n(3) xor C_BE_n(2) xor C_BE_n(1) xor C_BE_n(0);
end process PCI_Parity_Gen;

-- ***** �p���e�B�o�͐��� ***** --
PCI_Parity_Ctrl : process(PCICLK, RST_n)
begin
	if (RST_n = '0') then
		PAR_HiZ  <= '1';
		PAR_Port <= '0';
	elsif (PCICLK'event and PCICLK = '1') then
		if (PCIAD_HiZ = '0') then
			PAR_HiZ  <= '0';
			PAR_Port <= TGT_PAR;
		else
			PAR_HiZ  <= '1';
		end if;
		-- ��AD�o�X�̃h���C�u����1�N���b�N�x���PAR�𐧌�
	end if;
end process PCI_Parity_Ctrl;


end RTL;







